LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ConversorTemperatura IS
	PORT(
		xDados : IN STD_LOGIC_VECTOR  (7 DOWNTO 0);
		xTemp  : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END ConversorTemperatura;

ARCHITECTURE data_flow OF ConversorTemperatura IS

	SIGNAL RESULT_ONE : STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL RESULT_TWO : STD_LOGIC_VECTOR (15 DOWNTO 0);

BEGIN

	RESULT_ONE <= STD_LOGIC_VECTOR((UNSIGNED(xDados) * 10010110));
	RESULT_TWO <= STD_LOGIC_VECTOR((UNSIGNED(RESULT_ONE) / 11111111));
	
	xTemp      <= RESULT_TWO (15 DOWNTO 8);
	
END data_flow;